//###############################################
// Author:  Qazi Hamid Ullah (hamidullahqazi12@gmail.com)
// Date:    6/15/2023
// Module:  proc.v       
// Description: perform all operations
//  
//###############################################

module proc(DIN, Resetn, Clock, Run, DOUT, ADDR, W,r0);
    input [15:0] DIN;
    input Resetn, Clock, Run;
    output wire [15:0] DOUT;              //Data register 
    output wire [15:0] ADDR;              //address register
    output wire W;                        //it will enable both of write enable in memory and output reg enable
    output [15:0] r0;
    reg [15:0] BusWires;
    reg [3:0] Sel; // BusWires selector
    reg [0:7] Rin;  //enables of the register
    reg [15:0] Sum;
    reg IRin, ADDRin, Done, DOUTin, Ain, Gin, AddSub, ALUand;
    reg [2:0] Tstep_Q, Tstep_D;         //Tstep_Q present state and Tstep_D shows the next state
    wire [2:0] III, rX, rY; // instruction opcode and register operands
    wire [0:7] Xreg, Yreg;
    wire [15:0] R0, R1, R2, R3, R4, R5, R6, PC, A;      //A will hold one of the input to the ALU
    wire [15:0] G;          //it will hold the result of ALU
    wire [15:0] IR;         //Instr register 
    reg pc_inc, W_D;        
    wire IMM;               //it shows the 4th bit from right of the Instruction
    wire zero_flag, negative_flag;
	 reg carry_out_flag;          //for branch conditions
    reg carry_alu;         //carry out generated by ALU add/sub
    reg carr1;
	 wire out1, out2, out3;


    assign III = IR[15:13];
    assign IMM = IR[12];
    assign rX = IR[11:9];         //first register and also the destination register
    assign rY = IR[2:0];          //2nd register 
    //Enabling the specific registers enable signals according to instrcutions
    dec3to8 decX (rX, Xreg);
	 //dec3to8 decy (rX, Yreg);			//for branch instructions
	 
    parameter T0 = 3'b000, T1 = 3'b001, T2 = 3'b010, T3 = 3'b011, T4 = 3'b100, T5 = 3'b101;

    // Control FSM state table
    always @(Tstep_Q, Run, Done)          //Tstep_Q is present state and Tstep_D is next state 
        case (Tstep_Q)
            T0: // instruction fetch
                if (~Run) Tstep_D = T0;     //when run is 1 it will start
                else Tstep_D = T1;
            T1: // wait cycle for synchronous memory
                Tstep_D = T2;
            T2: // this time step stores the instruction word in IR
                Tstep_D = T3;
            T3: // some instructions end after this time step like mv or mvt  etc
                if (Done) Tstep_D = T0;
                else Tstep_D = T4;
            T4: // always go to T5 after this
                Tstep_D = T5;
            T5: // instructions end after this time step
                Tstep_D = T0;
            default: Tstep_D = 3'bxxx;
        endcase

    /* OPCODE format: III M XXX DDDDDDDDD, where 
    *     III = instruction, M = Immediate, XXX = rX. If M = 0, DDDDDDDDD = 000000YYY = rY
    *     If M = 1, DDDDDDDDD = #D is the immediate operand 
    *
    *  III M  Instruction   Description
    *  --- -  -----------   -----------
    *  000 0: mv   rX,rY    rX <- rY
    *  000 1: mv   rX,#D    rX <- D (0 extended)
    *  
    *  001 1: mvt  rX,#D    rX <- D << 8
    *  010 0: add  rX,rY    rX <- rX + rY
    *  010 1: add  rX,#D    rX <- rX + D
    *  011 0: sub  rX,rY    rX <- rX - rY
    *  011 1: sub  rX,#D    rX <- rX - D
    *  100 0: ld   rX,[rY]  rX <- [rY]
    *  101 0: st   rX,[rY]  [rY] <- rX
    *  110 0: and  rX,rY    rX <- rX & rY
    *  110 1: and  rX,#D    rX <- rX & D 
	 *  111 1: branch						*/
    parameter mv = 3'b000, mvt = 3'b001, add = 3'b010, sub = 3'b011, ld = 3'b100, st = 3'b101,
	     and_ = 3'b110, branch = 3'b111;
    // selectors for the BusWires multiplexer
    parameter Sel_R0 = 4'b0000, Sel_R1 = 4'b0001, Sel_R2 = 4'b0010, Sel_R3 = 4'b0011,
        Sel_R4 = 4'b0100, Sel_R5 = 4'b0101, Sel_R6 = 4'b0110, Sel_PC = 4'b0111, Sel_G = 4'b1000,
        Sel_D /* immediate data */ = 4'b1001, Sel_D8 /* immediate data << 8 */ = 4'b1010, 
        Sel_DIN /* data-in from memory */ = 4'b1011;
		parameter none = 3'b000, eq = 3'b001, ne = 3'b010, cc = 3'b011, cs = 3'b100, pl = 3'b101, mi = 3'b110;    //branch inst
		  
    // Control FSM outputs
    always @(*) begin
        // default values for control signals
        Done = 1'b0; Ain = 1'b0; Gin = 1'b0; AddSub = 1'b0; IRin = 1'b0; Sel = 4'bxxxx;
        DOUTin = 1'b0; ADDRin = 1'b0; W_D = 1'b0; Rin = 8'b0; pc_inc = 1'b0; ALUand = 1'b0;
        case (Tstep_Q)
            T0: begin // fetch the instruction
                Sel = Sel_PC; // put pc onto the internal bus
                ADDRin = 1'b1;
                pc_inc = Run; // to increment pc
            end
            T1: // wait cycle for synchronous memory
                ;
            T2: // store instruction on DIN in IR 
                IRin = 1'b1;
            T3: // define signals in T1
                case (III)
                    mv: begin
                        if (!IMM) Sel = rY;   // mv rX, rY
                        else Sel = Sel_D;     // mv rX, #D
                        Rin = Xreg;            //enable rX register
                        Done = 1'b1;
                    end
                    mvt: begin
                        // ... your code goes here
                        //here if the IMM bit is 1 mvt will proceed else wise branch instructions will process
     
                          Sel = Sel_D8;       //selecting the immediate value from MUX
                          Rin = Xreg;         //sending the enable signal of destination register
                          Done = 1'b1; end
                    branch: begin
                          //now branch instructions
                          //Sel = Sel_PC;
                          //Ain = 1'b1;
                         // if(IMM) begin
                          case(rX)
                            none:   Done = 1'b1;    //no branch 
                            eq:     if(zero_flag) begin    //it its true then insert the immediate address into PC
                                      Sel = Sel_D;     //insert the immediate data into buswires
                                      Rin[7] = 1'b1; 
                                      Done = 1'b1; end     //will enable PCin signal 
                                      else Done = 1'b1;
                            ne:      if(!zero_flag) begin
                                      Sel = Sel_D;
                                      Rin[7] = 1'b1;
                                      Done = 1'b1;  end 
                                      else Done = 1'b1; 
                            cc:      if(!carry_out_flag) begin
                                      Sel = Sel_D;
                                      Rin[7] = 1'b1;
                                      Done = 1'b1;  end
                                      else Done = 1'b1;
                            cs:      if(carry_out_flag) begin
                                      Sel = Sel_D;
                                      Rin[7] = 1'b1; 
                                      Done = 1'b1; end
                                      else Done = 1'b1;
                            pl:      if(!negative_flag) begin
                                      Sel = Sel_D;
                                      Rin[7] = 1'b1;  end
                            mi:      if(negative_flag) begin
                                      Sel = Sel_D;
                                      Rin[7] = 1'b1;  end       //pc enable*/
												  
                            default:  begin Sel = 4'bxxx; Rin = 8'd0; Done = 1'b0;end
                          endcase
                          //end
                          end
                    add, sub, and_: begin
                        // ... your code goes here
    //Here In this state we will select the RX register and save its value to Ain register
                        Sel = rX;     //rX register will be selected from MUX
                        Ain = 1'b1;   //rX data will go through bus to Ain
                    end
                    ld, st: begin
                        // ... your code goes here
    //load will load data from address RY to register RX
    //Store will save data from register RX to address RY
                        ADDRin = 1'b1;    //instruction will be read from memory RY address
                        Sel = rY;         //rY register content will be goto buswires 
                        //DOUTin = 1'b1;    //so that content at address rY move to Dout register
                    end
                    default:  begin 
						  Done = 1'b0; Ain = 1'b0; Gin = 1'b0; AddSub = 1'b0; IRin = 1'b0; Sel = 4'bxxxx;
						  DOUTin = 1'b0; ADDRin = 1'b0; W_D = 1'b0; Rin = 8'b0; pc_inc = 1'b0; ALUand = 1'b0;
						  end
                endcase
            T4: // define signals T2
                case (III)
                    add: begin
                        // ... your code goes here
                        Sel = (IMM) ? Sel_D : rY;     //if IMM = 1 then sel_D otherwise rY
                        Gin = 1'b1;                   //so that the ALU out can be stored in G

                    end
                    sub: begin
                        // ... your code goes here
                        Sel = (IMM) ? Sel_D : rY;     //if IMM = 1 then sel_D otherwise rY
                        AddSub = 1'b1;                //so that ALU can do subtraction
                        Gin = 1'b1;                   //so that the ALU out can be stored in G
                    end
                    and_: begin
                        // ... your code goes here
                        Sel = (IMM) ? Sel_D : rY;     //if IMM = 1 then sel_D otherwise rY
                        Gin = 1'b1;                   //so that the ALU out can be stored in G
                        ALUand = 1'b1;                //telling ALU to do AND
                    end
                    branch:  begin
                          //Sel = Sel_D8;
                          //Gin = 1'b1;
                          //Done = 1'b1;    
                    end


                    ld: // wait cycle for synchronous memory
                        ;
                    st: begin
                        // ... your code goes here
                        W_D = 1'b1;                   //so that data can be written in memory
                        Sel = rX;                     //so that data to be stord can be on Buswires
                        DOUTin = 1'b1;                //so that data can be written on memory
                        Done = 1'b1;
                    end
                    default:  begin Done = 1'b0; Ain = 1'b0; Gin = 1'b0; AddSub = 1'b0; IRin = 1'b0; Sel = 4'bxxxx;
        DOUTin = 1'b0; ADDRin = 1'b0; W_D = 1'b0; Rin = 8'b0; pc_inc = 1'b0; ALUand = 1'b0; end
                endcase
            T5: // define T3
                case (III)
                    add, sub, and_: begin
                        // ... your code goes here
                    //here we will write back the value of ALU into rX
                    Sel = Sel_G;     //will put ALU output into the Buswires
                    Rin = Xreg;     //will enable rX register
                    Done = 1'b1;     
                    end
                    ld: begin
                        // ... your code goes here
                        Rin = Xreg;       //will input the enable of RX-Destination register 
                        Done = 1'b1;
                        end
								 /*   branch:  begin
                          Sel = Sel_G;
                          Rin[7] = 1'b1;       //will enable PCin signal through the decoder
                          Done = 1'b1;
                    end*/
                    default:  begin Done = 1'b0; Ain = 1'b0; Gin = 1'b0; AddSub = 1'b0; IRin = 1'b0; Sel = 4'bxxxx;
        DOUTin = 1'b0; ADDRin = 1'b0; W_D = 1'b0; Rin = 8'b0; pc_inc = 1'b0; ALUand = 1'b0; end
                endcase
            default:  begin Done = 1'b0; Ain = 1'b0; Gin = 1'b0; AddSub = 1'b0; IRin = 1'b0; Sel = 4'bxxxx;
        DOUTin = 1'b0; ADDRin = 1'b0; W_D = 1'b0; Rin = 8'b0; pc_inc = 1'b0; ALUand = 1'b0; end
        endcase
    end   
   
    // Control FSM flip-flops
    always @(posedge Clock)
        if (!Resetn)
            Tstep_Q <= T0;
        else
            Tstep_Q <= Tstep_D;   
   
    regn reg_0 (BusWires, Rin[0], Clock, R0);
    regn reg_1 (BusWires, Rin[1], Clock, R1);
    regn reg_2 (BusWires, Rin[2], Clock, R2);
    regn reg_3 (BusWires, Rin[3], Clock, R3);
    regn reg_4 (BusWires, Rin[4], Clock, R4);
    regn reg_5 (BusWires, Rin[5], Clock, R5);
    regn reg_6 (BusWires, Rin[6], Clock, R6);
	 
    // R7 is program counter
    // module pc_count(R, Resetn, Clock, E, L, Q);
    pc_count pc (BusWires, Resetn, Clock, pc_inc, Rin[7], PC);

    regn reg_A (BusWires, Ain, Clock, A);
    regn reg_DOUT (BusWires, DOUTin, Clock, DOUT);
    regn reg_ADDR (BusWires, ADDRin, Clock, ADDR);
    regn reg_IR (DIN, IRin, Clock, IR);

    flipflop reg_W (W_D, Resetn, Clock, W);
    
    // alu
    always @(*)
        if (!ALUand)
            if (!AddSub)
                {carry_alu,Sum} = A + BusWires;
            else
                {carry_alu,Sum} = A - BusWires;
		  else
            Sum = A & BusWires;
    regn reg_G (Sum, Gin, Clock, G);

      //for carry out flag we must have registered carry_alu 
      always @ (posedge Clock) begin
        if(Gin)
          carry_out_flag <= carry_alu;
       // else 
         // carr1 <= 1'b0;   
      end
/*
    flipflop delay1 (carr1, Resetn, Clock, out1);
    flipflop delay2 (out1, Resetn, Clock, out2);
    flipflop delay3 (out2, Resetn, Clock, out3);
    flipflop delay4 (out3, Resetn, Clock, carry_out_flag);
      */
    //supporting the branch conditions beq, bneq etc 
      //creating flags for the branch conditions like zero flag, negative flag and carry out flag 
    
      assign zero_flag = (G == 0) ? 1 : 0;       //flag is 1 when ALU out put is 0
      assign negative_flag = (G[15]) ? 1 : 0;     //flag is 1 if the MSB (sign bit) is 1  
      //assign carry_out_flag = carry_alu;          //flag is 1 whenever carryout is generated in ALU the 



    // define the internal processor bus
    always @(*)
        case (Sel)
            Sel_R0: BusWires = R0;
            Sel_R1: BusWires = R1;
            Sel_R2: BusWires = R2;
            Sel_R3: BusWires = R3;
            Sel_R4: BusWires = R4;
            Sel_R5: BusWires = R5;
            Sel_R6: BusWires = R6;
            Sel_PC: BusWires = PC;
            Sel_G:  BusWires = G;
            Sel_D:  BusWires = {7'b0000000, IR[8:0]};
            Sel_D8: BusWires = {IR[7:0], 8'b00000000};
            default: BusWires = DIN;
        endcase


        assign r0 = R0;
endmodule



